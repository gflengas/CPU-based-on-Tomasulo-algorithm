library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Decoder5to32 is
    Port ( Awr : in  STD_LOGIC_VECTOR (4 downto 0);
           DecOut : out  STD_LOGIC_VECTOR (31 downto 0));
end Decoder5to32;

architecture Behavioral of Decoder5to32 is

begin
	process(Awr)
	begin
	case Awr is
	when "00000" => -- reg 0
		DecOut <= "00000000000000000000000000000000";
	
	when  "00001" => --reg 1 
		DecOut <= "00000000000000000000000000000010";
	
	when  "00010" => --reg 2
		DecOut <= "00000000000000000000000000000100";
	
	when  "00011" => --reg 3 
		DecOut <= "00000000000000000000000000001000";
	
	when  "00100" => --reg 4
		DecOut <= "00000000000000000000000000010000";
	
	when  "00101" => --reg 5
		DecOut <= "00000000000000000000000000100000";
	
	when  "00110" => --reg 6
		DecOut <= "00000000000000000000000001000000";
	
	when  "00111" => --reg 7 
		DecOut <= "00000000000000000000000010000000";
	
	when  "01000" => --reg 8
		DecOut <= "00000000000000000000000100000000";
	
	when  "01001" => --reg 9
		DecOut <= "00000000000000000000001000000000";
	
	when  "01010" => --reg 10
		DecOut <= "00000000000000000000010000000000";
		
	when  "01011" => --reg 11
		DecOut <= "00000000000000000000100000000000";

	when  "01100" => --reg 12
		DecOut <= "00000000000000000001000000000000";
	
	when  "01101" => --reg 13
		DecOut <= "00000000000000000010000000000000";
	
	when  "01110" => --reg 14
		DecOut <= "00000000000000000100000000000000";
	
	when  "01111" => --reg 15
		DecOut <= "00000000000000001000000000000000";
	
	when  "10000" => --reg 16
		DecOut <= "00000000000000010000000000000000";
	
	when  "10001" => --reg 17
		DecOut <= "00000000000000100000000000000000";
	
	when  "10010" => --reg 18
		DecOut <= "00000000000001000000000000000000";
	
	when  "10011" => --reg 19
		DecOut <= "00000000000010000000000000000000";
	
	when  "10100" => --reg 20
		DecOut <= "00000000000100000000000000000000";
	
	when  "10101" => --reg 21
		DecOut <= "00000000001000000000000000000000";
	
	when  "10110" => --reg 22
		DecOut <= "00000000010000000000000000000000";
	
	when  "10111" => --reg 23
		DecOut <= "00000000100000000000000000000000";
	
	when  "11000" => --reg 24
		DecOut <= "00000001000000000000000000000000";
	
	when  "11001" => --reg 25
		DecOut <= "00000010000000000000000000000000";
	
	when  "11010" => --reg 26
		DecOut <= "00000100000000000000000000000000";
	
	when  "11011" => --reg 27
		DecOut <= "00001000000000000000000000000000";
	
	when  "11100" => --reg 28
		DecOut <= "00010000000000000000000000000000";
	
	when  "11101" => --reg 29
		DecOut <= "00100000000000000000000000000000";
	
	when  "11110" => --reg 30
		DecOut <= "01000000000000000000000000000000";
	
	when  others => --reg 31
		DecOut <= "10000000000000000000000000000000";
	
	end case;
	
	end process ;
end Behavioral;

